module timer #(parameter WAIT_TIME = 434) (
	input clk, rst,
	output reg done
);

int WIDTH = $clog2(WAIT_TIME),
reg [WIDTH-1 : 0] counter;
	
always_ff @(posedge clk) begin
	if (rst) begin
		counter <= '0;
		done <= 1'b0;
	end
	else if (counter < WAIT_TIME)
		counter <= counter + 1'b1;
	else begin
		counter <= '0;
		done <= 1'b1;
	end

end
endmodule
